module Syncrhonizer(input logic clock, input logic reset, input logic resetButton,
                    input logic recordButton, input logic playButton, input logic clipRecordNum,
                    input logic clipPlayNum, output logic resetBSync, output logic recordBSync,
                    output logic playBSync, output logic clipRSync, output logic clipPSync);

endmodule
