module Timer(input logic clock, input logic reset, input logic isEnabled, output logic secondMarker);

endmodule
