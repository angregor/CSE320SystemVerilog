module LEDinterface(input logic clock, input logic reset, input logic clipNum, input logic recordOrPlay,
                    output logic[6:0] cathode, output logic A0, output logic A7);

endmodule
