module Controller(input logic clock, input logic reset, input logic resetButtonS,
                    input logic recordButtonS, input logic playButtonS, input logic clipRecordNumS,
                    input logic clipPlayNumS, output logic resetBSync, output logic isEnabledTimer,
                    output logic enableDeSerial, output logic enableSerial, output memAddress);

endmodule
