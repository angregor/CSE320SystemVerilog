module clockScalar(input logic clock, input logic reset, output logic scaledClock);

endmodule
