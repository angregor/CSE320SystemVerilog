module addressCounter(input logic clock, input logic reset, input logic desDone, input logic sDone,
                      output logic[15:0] address);

endmodule
