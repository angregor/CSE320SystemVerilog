module Syncrhonizer(input logic clock, input logic reset, input logic resetButton, input logic clipNum, input logic playOrRecord, input logic ActionButton,
  output logic ActionSync, output logic ClipNumSync, output logic PlayOrRecordSync, output logic resetButtonSync);

endmodule
